library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ROM is
	Generic (
		N : positive := 6;		--address length
		M : positive := 32);	--data word length
	Port (
		ADDR     :  in STD_LOGIC_VECTOR (N-1 downto 0);
		DATA_OUT : out STD_LOGIC_VECTOR (M-1 downto 0));
end ROM;

architecture Behavioral of ROM is

type ROM_array is array (0 to 2**N-1) of STD_LOGIC_VECTOR (M-1 downto 0);

constant ROM : ROM_array := (
	X"E2C00000", X"E2801005", X"E1E02001", X"E0513002",	-- 1h 16ada
	X"0A000000", X"51814003", X"E0015004", X"E5801004",
	X"EB00000F", X"E1A0A089", X"E1A000A0", X"E5906004",
	X"E2267009", X"E357000D", X"B2808050", X"E5808024",
	
	X"E08FF000", X"E3E02000", X"E590F024", X"EAFFFFEB",	-- 2h 16ada
	X"E245B00A", X"E28BC007", X"E1A0DFEC", X"E0C00000",
	X"EAFFFFE6", X"E2800001", X"E1B09141", X"62800064",
	X"22405032", X"E0C0F00E", X"00000000", X"00000000",
	
	X"00000000", X"00000000", X"00000000", X"00000000",	-- 3h 16ada
	X"00000000", X"00000000", X"00000000", X"00000000",
	X"00000000", X"00000000", X"00000000", X"00000000",
	X"00000000", X"00000000", X"00000000", X"00000000",
	
	X"00000000", X"00000000", X"00000000", X"00000000",	-- 4h 16ada
	X"00000000", X"00000000", X"00000000", X"00000000",
	X"00000000", X"00000000", X"00000000", X"00000000",
	X"00000000", X"00000000", X"00000000", X"00000000"
	);

begin

	DATA_OUT <= ROM(to_integer(unsigned(ADDR)));

end Behavioral;